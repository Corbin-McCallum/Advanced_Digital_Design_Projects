library ieee;
use ieee.std_logic_1164.all;

entity top_level is
	
end entity top_level;

architecture arch1 of top_level is

begin

end architecture top_level;